-- Criando um somador de quatro bits com quatro somadores de um bit usando port map
