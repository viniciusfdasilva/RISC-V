library ieee;
use ieee.std_logic_1164.all;

entity alu is
	port(
		inputA : in std_logic;
		inputB : in std_logic;
		output : out std_logic
	);
end alu;

architecture alu of alu is
begin
end alu;